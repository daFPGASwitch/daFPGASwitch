module top #()
(
    // egress
); 



// pack_gen(0)
// pack_gen(1)
// pack_gen(2)
// pack_gen(3)


