// Inside of egress

module pack_val #()
(
    input meta
)

endmodule